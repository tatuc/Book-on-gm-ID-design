** sch_path: /foss/designs/Book-on-gm-ID-design/starter_files_open_source_tools/ihp-sg13g2/techsweep_sg13_hv_nmos.sch
**.subckt techsweep_sg13_hv_nmos
vg g 0 DC 0.6 AC 1
vd d 0 1.65
vb b 0 0
Hn n 0 vd 1
XM1 d g 0 b sg13_hv_nmos w={wx} l={lx} ng=1 m=1
**** begin user architecture code


.param wx=5u lx=0.35u
.op

.control
option numdgt = 3
set wr_singlescale
set wr_vecnames

compose l_vec  values 0.45u 0.5u 0.55u
+ 0.6u 0.7u 0.8u 0.9u 1u 2u 3u
compose vg_vec start= 0 stop=3.301  step=25m
compose vd_vec start= 0 stop=3.301  step=25m
compose vb_vec start= 0 stop=-0.6   step=-0.2

foreach var1 $&l_vec
  alterparam lx=$var1
  reset
  foreach var2 $&vg_vec
    alter vg $var2
    foreach var3 $&vd_vec
      alter vd $var3
      foreach var4 $&vb_vec
        alter vb $var4
        run
        wrdata techsweep_sg13_hv_nmos.txt all
        destroy all
        set appendwrite
        unset set wr_vecnames
      end
    end
  end
end
unset appendwrite

alterparam lx=0.35u
reset
op
show
write techsweep_sg13_hv_nmos.raw
.endc




.save @n.xm1.nsg13_hv_nmos[cdd]
.save @n.xm1.nsg13_hv_nmos[cgb]
.save @n.xm1.nsg13_hv_nmos[cgd]
.save @n.xm1.nsg13_hv_nmos[cgdol]
.save @n.xm1.nsg13_hv_nmos[cgg]
.save @n.xm1.nsg13_hv_nmos[cgs]
.save @n.xm1.nsg13_hv_nmos[cgsol]
.save @n.xm1.nsg13_hv_nmos[cjd]
.save @n.xm1.nsg13_hv_nmos[cjs]
.save @n.xm1.nsg13_hv_nmos[css]
.save @n.xm1.nsg13_hv_nmos[gds]
.save @n.xm1.nsg13_hv_nmos[gm]
.save @n.xm1.nsg13_hv_nmos[gmb]
.save @n.xm1.nsg13_hv_nmos[ids]
.save @n.xm1.nsg13_hv_nmos[l]
.save @n.xm1.nsg13_hv_nmos[sfl]
.save @n.xm1.nsg13_hv_nmos[sid]
.save @n.xm1.nsg13_hv_nmos[vth]
.save @vb[dc]
.save @vd[dc]
.save @vg[dc]
.save g d b n


 .lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt
**** end user architecture code
**.ends
.end
